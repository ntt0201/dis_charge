** circuit: digital_BGR_model
** -------- discharge network description -------- **
.subckt discharge_nwk ctrl _VP_ VGND W=0.5
XM1 net3 net3 _VP_ _VP_ sky130_fd_pr__pfet_01v8 L=0.15 W="W" nf=1
XM2 net2 net2 net1 net1 sky130_fd_pr__pfet_01v8 L=0.15 W="W" nf=1
XM3 net1 net1 net3 net3 sky130_fd_pr__pfet_01v8 L=0.15 W="W" nf=1 
XM4 net4 net4 net2 net2 sky130_fd_pr__pfet_01v8 L=0.15 W="W" nf=1
XM5 netk netk net4 net4 sky130_fd_pr__pfet_01v8 L=0.15 W="W" nf=1
XC1 _VP_ VGND sky130_fd_pr__cap_mim_m3_2 W=14.5 L=1.5 MF=10 m=10
XMk netk ctrl VGND VGND sky130_fd_pr__nfet_01v8 L=0.15 W=2 nf=2
.ends
X_discharge_nwk ctrl VP GND discharge_nwk W=W
*charge sw 
asw a_charge_sw %gd(VP_ VP) switch3
.model switch3 aswitch(cntl_off='v_dd/2-5m' cntl_on='v_dd/2+5m' r_off=1e15
+ r_on=10k log=TRUE limit=TRUE)
** -------- end discharge network description --------**

** -------- Time to digital description ---------- **
X_counter1 d_clk d_low d_rst o0 o1 o2 o3 o4 o5 o6 o7 o8 o9 o10 o11 o12 o13 o14 o15 counter_16b
ECMP a_fb_cmp net3 TABLE {V(ref_sig ,VP)} = ( -1mV , 0V ) ( 1mV , 0.8V )
r1 VDD ref_sig 30k
r2 ref_sig gnd 10k
r3 net3 gnd 10k
** -------- end 

** ---------------- DAC description --------------- **

V_DAC VP_ gnd DC = 0.05
* r5 r_in_dac gnd 1k 
** ----------------- end

** ---------- Simulation controller description ----------- **

X_rst d_clk d_low d_rst0 d_fb_cmp d_rst d_rst_bar bit9 bit10 set_dac_sig d_charge_sw bit_sel0 bit_sel1 controller

.subckt controller clk low rst0 cmp_sig rst rst_bar bit9 bit10 set_dac_sig charge_sw bit_sel0 bit_sel1
a_or0 [rst0 rst1] rst or1
a_dff0 d0 cmp_sig low rst0 sig1 d0 flop1
a_dff1 d1 bit11 low rst0 sig2 d1 flop1
a_xor0 [sig1 sig2] rst1 xor1
a_inv0 rst1 rst1_bar inv1
a_inv1 rst1_bar rst1_dl inv1

X_counter2 clk low rst1_bar bit8 bit9 bit10 bit11 counter_12b
a_and0 [bit8 ~bit9 ~bit10] set_dac_sig and1
a_and1 [~bit11 bit10] charge_sw2 and1
a_or1 [rst0 charge_sw2] charge_sw or1
x_sub_cnt rst low rst0 bit_sel0 bit_sel1 counter_2b

.model and1 d_and(rise_delay = 0.5e-9 fall_delay = 0.3e-9 input_load = 0.5e-12)
.model inv1 d_inverter(rise_delay = 0.5e-9 fall_delay = 0.3e-9 input_load = 0.5e-12)
.model or1 d_or(rise_delay = 0.5e-9 fall_delay = 0.3e-9 input_load = 0.5e-12)
.model flop1 d_dff(clk_delay = 13.0e-9 set_delay = 25.0e-9 reset_delay = 27.0e-9 
+ ic = 2 rise_delay = 10.0e-9 fall_delay = 3e-9)
.model nand1 d_nand(rise_delay = 0.5e-9 fall_delay = 0.3e-9 input_load = 0.5e-12)
.model xor1 d_xor(rise_delay = 0.5e-9 fall_delay = 0.3e-9 input_load = 0.5e-12)
.ends

abridge1 [d_charge_sw] [a_charge_sw] dac1
.model dac1 dac_bridge(out_low = 0 out_high = 'v_dd' out_undef = 'v_dd/2'
+ input_load = 5.0e-12 t_rise = 0.5e-9
+ t_fall = 0.5e-9)

*** adc_bridge blocks ***
aconverter [a_clk  a_rst0 a_fb_cmp a_high a_sig 0] [d_clk d_rst0 d_fb_cmp d_hi d_sig d_low] adc1
.model adc1 adc_bridge (in_low='v_dd/2-5m' in_high='v_dd/2+5m' rise_delay=1.0e-12 fall_delay=1.0e-12)

* Voltage setup for the circuit
V_sup VDD GND DC = 'v_dd'
V_clk a_clk GND pulse (0 'v_dd' 0 'prd/20' 'prd/20' '9*prd/20' prd)
V_rst0 a_rst0 net4 pulse  (0 'v_dd' 'T_set' 1e-12 1e-12 'T_on' 1 1)
r4 net4 gnd 10k
V_ctrl ctrl net6 dc = 'v_dd'
r6 net6 gnd 10k 
*input sources resistance

* Setup simulation 
*.lib ~/work/conda_eda/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.lib /home/dkits/efabless/mpw-7a/pdks/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.inc ./../lib/counter.spice
.inc ./../lib/mux2i_1.spice
.param clk_freq = 0.5e6
.param prd = '1/clk_freq'
.param T_set = 0.22m T_on = 0.5m
.param W = 0.5
.param V_init = 0.2
.param v_dd = 0.555
.csparam v_dd_ = {v_dd}
.ic v(VP) = V_init
.option trtol = 5
.save vp vp_ a_rst0 a_charge_sw x_rst.bit_sel0 x_rst.bit_sel1 d_rst set_dac_sig
+ ctrl
+ o15 o14 o13 o12 o11 o10 o9 o8 o7 o6 o5 o4 o3 o2 o1 o0
.temp 29
** -------------------- end controller descriptions ----------------------- **
.control
echo  ______________________________________
echo |   go to the measurement operation    |
echo  --------------------------------------
let NoL = 4096			$ Number of DAC Levels
let m = vector(3)		$ storage of DAC m levels
let n = vector(3)		$ storage of TDC discharge time
let DAC_vol = vector(3)		$ storage of the DAC voltage

* get the value of the m vector
let ix = 0
while (ix<3)
	let m[ix] = `/bin/bash -c "python processor_model.py $&ix"`
	let DAC_vol[ix] = (m[ix]/NoL)*v_dd_
	let ix = ix+1
end

let half_vdd = v_dd_/2
stop when v(a_rst0)>'$&half_vdd'  when v(VP_)<0.1
let cnt_stop=1
let dvol1 = DAC_vol[0]-0.01
stop when set_dac_sig=1  when bit_sel0=0 when bit_sel1=0 when v(VP_)>'$&dvol1'
let dvol2 = DAC_vol[1]-0.01
stop when set_dac_sig=1  when bit_sel0=1 when bit_sel1=0 when v(VP_)>'$&dvol2'
stop when set_dac_sig=1  when bit_sel0=0 when bit_sel1=1 when v(ctrl)>'$&half_vdd'

tran 100n 75m

alter V_DAC dc = dac_vol[0]
resume
eprint o15 o14 o13 o12 o11 o10 o9 o8 o7 o6 o5 o4 o3 o2 o1 o0 > stop1.txt
alter V_DAC dc = dac_vol[1]
resume
eprint o15 o14 o13 o12 o11 o10 o9 o8 o7 o6 o5 o4 o3 o2 o1 o0 > stop2.txt
alter V_DAC dc = dac_vol[2]
resume
eprint o15 o14 o13 o12 o11 o10 o9 o8 o7 o6 o5 o4 o3 o2 o1 o0 > stop3.txt
let m_ref = `/bin/bash -c "python processor_model.py 3"`
let DAC_ref = (m_ref/NoL)*v_dd_
alter V_DAC dc = dac_ref
alter V_ctrl dc = 0 
resume
plot VP VP_ d_rst
.endc
.GLOBAL GND
.end

