** circuit: digital_BGR_model

.subckt discharge_nwk VP VGND 
XM1 net3 net3 VP VP sky130_fd_pr__pfet_01v8 L=0.15 W="W" nf=1
XM2 net2 net2 net1 net1 sky130_fd_pr__pfet_01v8 L=0.15 W="W" nf=1
XM3 net1 net1 net3 net3 sky130_fd_pr__pfet_01v8 L=0.15 W="W" nf=1 
XM4 net4 net4 net2 net2 sky130_fd_pr__pfet_01v8 L=0.15 W="W" nf=1
XM5 GND VGND net4 net4 sky130_fd_pr__pfet_01v8 L=0.15 W="W" nf=1
XC1 VP VGND sky130_fd_pr__cap_mim_m3_2 W=14.5 L=1.5 MF=10 m=10
.ends
 
* Digital circuits by xspice
a8 enb %gd(VP_ VP) switch3

.model switch3 aswitch(cntl_off=0.0 cntl_on=0.4 r_off=1e15
+ r_on=10k log=TRUE limit=TRUE)


* Voltage setup for the circuit
V_DAC VP_ GND DC=0.8
V_sup VDD GND DC=0.8
V_enb enb GND pulse (0 V_on T_set 0 0 T_on 40m 1)
V_clk clk GND pulse (0 0.8 0 'prd/20' 'prd/20' '9*prd/20' prd)

* Setup simulation 
.lib ~/work/conda_eda/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.param clk_freq = 1e6
.param prd = '1/clk_freq'
.param T_set = 0.1m T_on = 1m V_on = 0.4
.param W = 0.5
.param V_init = 0.2
.ic v(VP) = V_init

.tran 100n 40m

.control
save VP_ VP enb clk  
set N = 65536
let DAC_vol = ($m_set/$N)*$v_dd
alter V_sup dc=$v_dd
alter V_DAC dc=DAC_vol
run
let ix=ix+1
meas tran DAC_out AVG v(VP_) from=2m to=10m
print DAC_out
end
	write d_bgr_model.raw
else
	echo "go to the meas op"
	let m = vector(3)
	let n = vector(3)
	let m[0] = $m1
	let m[1] = $m2
	let m[2] = $m3
	let im = 0
	while im<3
	  let DAC_vol = (m[im]/$N)*$v_dd
	  alter V_DAC dc=DAC_vol
	  alter V_sup dc=$v_dd
	  run
	  let quad_dd = $v_dd/4
	  meas tran DAC_out AVG v(VP_) from=2m to=10m
	  meas tran t_dis WHEN v(VP)=quad_dd CROSS=LAST
	*  meas tran t_dis trig v(enb) val=0 FALL=1  targ v(VP) val=quad_dd FALL=1
	  let n[im] = 't_dis-1.1m'
	  print DAC_out
	  let im = im+1
	end
	print n > discharge_time.txt
	write d_bgr_model.raw
end
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
